package eth_tb_pkg;
  import uvm_pkg::*;
  `include "eth_tb_scoreboard.sv"
  `include "eth_tb_vsequencer.sv"
  `include "eth_tb_vseq.sv"
  `include "eth_tb.sv"
endpackage

`include "tc_basic.sv"

package apb_pkg;
  import uvm_pkg::*;
  `include "apb_trans.sv"
endpackage

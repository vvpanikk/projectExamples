package eth_pkg;
  import uvm_pkg::*;
  `include "eth_trans.sv"
  `include "eth_config.sv"
  `include "eth_sequencer.sv"
  `include "eth_driver.sv"
  `include "eth_monitor.sv"
  `include "eth_agent.sv"
  `include "eth_env.sv"
  `include "eth_seq.sv"
endpackage
